/*
 * Verilog module for 32-Bit ALU based on SPARC Architecture.
 * Written by Johnny Sanchez - Github username:johnnyrsm
 */
module ALU(output reg [31:0] Out, output reg C, N, V, Z, input [31:0] A, B, input [5:0] OpCode, input Cin);

//*************************************
//	OpCode definitions
//	for each Instruction
//*************************************

//*************************************
//	Basic Arithmetic
//	Instructions
//*************************************

parameter [5:0] ADD = 6'b000000,
		ADDCC = 6'b010000,
		ADDX = 6'b001000,	
		ADDXCC = 6'b011000,
		SUB = 6'b000100,
		SUBCC = 6'b010100,
		SUBX = 6'b001100,
		SUBXCC = 6'b011100,

//************************************
//	Logical
//	Instructions
//************************************

		AND = 6'b000001,
		ANDCC = 6'b010001,
		ANDN = 6'b000101,
		ANDNCC = 6'b010101,	
		OR = 6'b000010,		
		ORCC = 6'b010010,
		ORN = 6'b000110,
		ORNCC = 6'b010110,
                XOR = 6'b000011,
                XORCC = 6'b010011,
                XORN = 6'b000111,
                XORNCC = 6'b010111,

//************************************
//	Shift Instructions
//************************************

		SLL = 6'b100101,	
		SRL = 6'b100110,	
		SRA = 6'b100111,

//***********************************
//	Load/Store
//	Instructions
//***********************************

		LSB = 6'b001001,
		LDSH = 6'b001010,
		LD = 6'b001000,
		LDUB = 6'b000001,
		LDUH = 6'b000010,
		LDD = 6'b000011,
		STB = 6'b000101,
		STH = 6'b000110,
		ST = 6'b000100,
		STD = 6'b000111;

always@(OpCode, A, B)
begin
        case(OpCode)
//-----------------------------------
//---Basic-Arithmetic-Instructions---
//-----------------------------------

        ADD:
        begin
                Out = A + B;
        end

        ADDCC:
        begin
                Out = A + B;
                N = Out[31];

                if(A + B > 32'hFFFFFFFF)
                        C = 1'b1;
                else
                        C = 1'b0;

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;

                if((A[31] == B[31]) && (A[31] != Out[31]))
                        V = 1'b1;
                else
                        V = 1'b0;
	end

	ADDX:
	begin
		Out = A + B + Cin;
	end
	
	ADDXCC:
	begin
		Out = A + B + Cin;
                N = Out[31];

                if(A + B + Cin > 32'hFFFFFFFF)
                        C = 1'b1;
                else
                        C = 1'b0;

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;

                if((A[31] == B[31]) && (A[31] != Out[31]))
                        V = 1'b1;
                else
                        V = 1'b0;
	end

	SUB:
	begin
		Out = A - B;
	end

	SUBCC:
	begin
		Out = A - B;
		N = Out[31];

		if(B > A)
                        C = 1'b1;
                else
                        C = 1'b0;

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;

                if((A[31] != B[31]) && (A[31] != Out[31]))
                        V = 1'b1;
                else
                        V = 1'b0;

	end
	
	SUBX:
	begin
		Out = A - B - Cin;
	end

	SUBXCC:
	begin
		Out = A - B - Cin;
		N = Out[31];

                if(B > A)
                        C = 1'b1;
                else
                        C = 1'b0;

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;

                if((A[31] != B[31]) && (A[31] != Out[31]))
                        V = 1'b1;
                else
                        V = 1'b0;

	end

//-----------------------------
//---Logical-Instructions------
//-----------------------------
	
	AND:
	begin
		Out = A & B;
	end

	ANDCC:
	begin
		Out = A & B;
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
		
		C = ~Z;
		V = 0;
		
	end
	
	ANDN:
	begin
		Out = A & (~B);
	end

	ANDNCC:
	begin
		Out = A & (~B);
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
		
		C = ~Z;
		V = 0;
		
	end
	
	OR:
	begin
		Out = A | B;
	end

	ORCC:
	begin
		Out = A | B;
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
               
                C = ~Z;
                V = 0;
              
	end

	ORN:
	begin
		Out = A | (~B); 
	end

	ORNCC:
	begin
		Out = A | (~B);
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
               
                C = ~Z;
                V = 0;
                
	end

	XOR:
	begin
		Out = A ^ B; 
	end
	
	XORCC:
	begin
		Out = A ^ B;
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
                
                C = ~Z;
                V = 0;
                
	end

	XORN:
	begin
		Out = A ^ (~B);
	end

	XORNCC:
	begin
		Out = A ^ (~B);
		N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
                
                C = ~Z;
                V = 0;
                
	end

//--------------------------
//---Shift-Instructions-----
//--------------------------

	SLL:
	begin
		Out = A << (B & 32'h0000001F);
                N = Out[31];
 
                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
                 
                C = ~Z;
                V = 0;  
	end
		
	SRL:
	begin
		Out = A >> (B & 32'h0000001F);
                N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
                
                C = ~Z;
                V = 0;  
	end

	SRA:
	begin
		Out = A >>> (B & 32'h0000001F);
                N = Out[31];

                if(Out == 0)
                        Z = 1'b1;
                else
                        Z = 1'b0;
                 
                C = ~Z;
                V = 0;  
	end

//------------------------------
//---Load/Store-Instructions----
//------------------------------

/*
 * Load instructions produce an Effective
 * Address from the sum of its operands
 */
	LSB:
	begin
		Out = A + B;		
	end

	LDSH:
	begin
		Out = A + B;
	end

	LD:
	begin
		Out = A + B;
	end

	LDUB:
	begin
		Out = A + B;
	end

	LDUH:
	begin
		Out = A + B;
	end

	LDD:
	begin
		Out = A + B;
	end

/*
 * Store instructions produce an Effective
 * Address from the sum of its operands
 */
	STB:
	begin
		Out = A + B;
	end

	STH:
	begin
		Out = A + B;
	end
	
	ST:
	begin
		Out = A + B;
	end

	STD:
	begin
		Out = A + B;
	end

end
endmodule
